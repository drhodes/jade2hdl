------------------------------------------------------------------
-- VHDL PRELUDE --------------------------------------------------

-- library IEEE;
-- use IEEE.STD_LOGIC_1164.ALL;

-- entity mod_user_and2 is
--   port (a : in std_logic_vector(0 downto 0);
--         b : in std_logic_vector(0 downto 0);
--         vout : out std_logic_vector(0 downto 0));
-- end entity mod_user_and2 ;
-- architecture behavioral of mod_user_and2 is
-- begin
--     vout <= a and b;
-- end architecture behavioral ;

-- /gates/and4 ------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity mod_gates_and4 is
  port (a : in std_logic_vector(0 downto 0);
        b : in std_logic_vector(0 downto 0);
        c : in std_logic_vector(0 downto 0);
        d : in std_logic_vector(0 downto 0);
        vout : out std_logic_vector(0 downto 0));
end entity mod_gates_and4 ;
architecture behavioral of mod_gates_and4 is
begin
  vout <= a and b and c and d;
end architecture behavioral ;

-- /gates/and2 ------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity mod_gates_and2 is
  port (a : in std_logic_vector(0 downto 0);
        b : in std_logic_vector(0 downto 0);
        vout : out std_logic_vector(0 downto 0)) ;
end entity mod_gates_and2 ;
architecture behavioral of mod_gates_and2 is
begin
  vout <= a and b;
end architecture behavioral ;

-- /gates/buffer ------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity mod_gates_buffer is
  port (a : in std_logic_vector(0 downto 0);
        vout : out std_logic_vector(0 downto 0)) ;
end entity mod_gates_buffer ;
architecture behavioral of mod_gates_buffer is
begin
  vout <= a;
end architecture behavioral ;


-- /gates/or2 ------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity mod_gates_or2 is
  port (a : in std_logic_vector(0 downto 0);
        b : in std_logic_vector(0 downto 0);
        vout : out std_logic_vector(0 downto 0)) ;
end entity mod_gates_or2 ;
architecture behavioral of mod_gates_or2 is
begin
  vout <= a or b;
end architecture behavioral ;


-- END VHDL PRELUDE ----------------------------------------------
------------------------------------------------------------------
